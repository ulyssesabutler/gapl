//
// Copyright (C) 2019 Yuta Tokusashi
// All rights reserved.
//
// This software was developed by
// Stanford University and the University of Cambridge Computer Laboratory
// under National Science Foundation under Grant No. CNS-0855268,
// the University of Cambridge Computer Laboratory under EPSRC INTERNET Project EP/H040536/1 and
// by the University of Cambridge Computer Laboratory under DARPA/AFRL contract FA8750-11-C-0249 ("MRC2"), 
// as part of the DARPA MRC research programme.
//
// @NETFPGA_LICENSE_HEADER_START@
//
// Licensed to NetFPGA C.I.C. (NetFPGA) under one or more contributor
// license agreements.  See the NOTICE file distributed with this work for
// additional information regarding copyright ownership.  NetFPGA licenses this
// file to you under the NetFPGA Hardware-Software License, Version 1.0 (the
// "License"); you may not use this file except in compliance with the
// License.  You may obtain a copy of the License at:
//
//   http://www.netfpga-cic.org
//
// Unless required by applicable law or agreed to in writing, Work distributed
// under the License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied.  See the License for the
// specific language governing permissions and limitations under the License.
//
// @NETFPGA_LICENSE_HEADER_END@
//

// This file is generated by ./gen.sh
module ncams #(
	parameter MEM_TYPE         = 1,
	parameter CAM_MODE         = 0,
	parameter ID_BITS          = 1,
    parameter TCAM_ADDR_WIDTH  = 5 ,
    parameter TCAM_DATA_WIDTH  = 32,
    parameter TCAM_ADDR_TYPE   = 0,
    parameter TCAM_MATCH_ADDR_WIDTH = 5
)(
	input  wire                       	    clk,
	input  wire                       	    rst,
    input  wire                             we,
    input  wire [TCAM_ADDR_WIDTH+ID_BITS-1:0]       addr_wr,
    input  wire [TCAM_DATA_WIDTH-1:0]       din,
    output wire                             busy,
    input  wire [TCAM_DATA_WIDTH-1:0]       cmp_din,
    output wire                             match,
    output wire [TCAM_MATCH_ADDR_WIDTH+ID_BITS-1:0] match_addr
);

/* 
 * wires 
 */

 (* dont_touch="true" *) reg                             we_0;
 (* dont_touch="true" *) reg [TCAM_ADDR_WIDTH+ID_BITS-1:0]       addr_wr_0;
 (* dont_touch="true" *) reg [TCAM_DATA_WIDTH-1:0] 	     din_0;
 (* dont_touch="true" *) reg [TCAM_DATA_WIDTH-1:0] 	     cmp_din_0;
 (* dont_touch="true" *) wire                       	     busy_0;
 (* dont_touch="true" *) wire 				             match_0;
 (* dont_touch="true" *) wire [TCAM_MATCH_ADDR_WIDTH-1:0] match_addr_0;

 (* dont_touch="true" *) reg                             we_1;
 (* dont_touch="true" *) reg [TCAM_ADDR_WIDTH+ID_BITS-1:0]       addr_wr_1;
 (* dont_touch="true" *) reg [TCAM_DATA_WIDTH-1:0] 	     din_1;
 (* dont_touch="true" *) reg [TCAM_DATA_WIDTH-1:0] 	     cmp_din_1;
 (* dont_touch="true" *) wire                       	     busy_1;
 (* dont_touch="true" *) wire 				             match_1;
 (* dont_touch="true" *) wire [TCAM_MATCH_ADDR_WIDTH-1:0] match_addr_1;

reg [3:0] rst_vct;
always @ (posedge clk) begin
	rst_vct <= rst ? 4'b1111 : 4'b0000;
end

always @ (posedge clk) 
	if (!rst_vct[0]) begin
		we_0 <= 0;
		addr_wr_0 <= 0;
		din_0 <= 0;
		cmp_din_0 <= 0;
	end else begin
		we_0 <=  we ;
		addr_wr_0 <=  addr_wr ;
		din_0 <= din;
		cmp_din_0 <= cmp_din;
	end

always @ (posedge clk) 
	if (!rst_vct[1]) begin
		we_1 <= 0;
		addr_wr_1 <= 0;
		din_1 <= 0;
		cmp_din_1 <= 0;
	end else begin
		we_1 <=  we ;
		addr_wr_1 <=  addr_wr ;
		din_1 <= din;
		cmp_din_1 <= cmp_din;
	end


assign busy = busy_0 & busy_1;

/*
 * CAM instances
 */
(* keep_hierarchy="yes" *) cam_w #(
	.ID                       (0),
	.ID_BITS                  (ID_BITS),
	.MEM_TYPE                 (MEM_TYPE),
	.CAM_MODE                 (CAM_MODE),
	.C_TCAM_ADDR_WIDTH  	  (TCAM_ADDR_WIDTH), 
	.C_TCAM_DATA_WIDTH   	  (TCAM_DATA_WIDTH), 
	.C_TCAM_ADDR_TYPE	      (TCAM_ADDR_TYPE),
	.C_TCAM_MATCH_ADDR_WIDTH  (TCAM_MATCH_ADDR_WIDTH)
) u_cam_0 (
	.CLK         (clk),             //input					
	.WE          ((addr_wr_0[ID_BITS-1:0] == 0)?we_0:0),         //input					
	.ADDR_WR     ((addr_wr_0[ID_BITS-1:0] == 0)?addr_wr_0[ID_BITS+TCAM_ADDR_WIDTH-1:ID_BITS]:0),    //input   [C_TCAM_ADDR_WIDTH-1:0]	
	.DIN         (din_0),        //input   [C_TCAM_DATA_WIDTH-1:0]	
	.BUSY        (busy_0),       //output        			

	.CMP_DIN     (cmp_din_0),    //input   [C_TCAM_DATA_WIDTH-1:0]	
	.MATCH       (match_0),      //output         			
	.MATCH_ADDR  (match_addr_0)  //output  [C_TCAM_MATCH_ADDR_WIDTH-1:0]	
);

(* keep_hierarchy="yes" *) cam_w #(
	.ID                       (1),
	.ID_BITS                  (ID_BITS),
	.MEM_TYPE                 (MEM_TYPE),
	.CAM_MODE                 (CAM_MODE),
	.C_TCAM_ADDR_WIDTH  	  (TCAM_ADDR_WIDTH), 
	.C_TCAM_DATA_WIDTH   	  (TCAM_DATA_WIDTH), 
	.C_TCAM_ADDR_TYPE	      (TCAM_ADDR_TYPE),
	.C_TCAM_MATCH_ADDR_WIDTH  (TCAM_MATCH_ADDR_WIDTH)
) u_cam_1 (
	.CLK         (clk),             //input					
	.WE          ((addr_wr_1[ID_BITS-1:0] == 1)?we_1:0),         //input					
	.ADDR_WR     ((addr_wr_1[ID_BITS-1:0] == 1)?addr_wr_1[ID_BITS+TCAM_ADDR_WIDTH-1:ID_BITS]:0),    //input   [C_TCAM_ADDR_WIDTH-1:0]	
	.DIN         (din_1),        //input   [C_TCAM_DATA_WIDTH-1:0]	
	.BUSY        (busy_1),       //output        			

	.CMP_DIN     (cmp_din_1),    //input   [C_TCAM_DATA_WIDTH-1:0]	
	.MATCH       (match_1),      //output         			
	.MATCH_ADDR  (match_addr_1)  //output  [C_TCAM_MATCH_ADDR_WIDTH-1:0]	
);

/*
 * Priority Encoder instances
 */

(* dont_touch="true" *) wire [TCAM_MATCH_ADDR_WIDTH+ID_BITS-1:0] l1_prio_match_addr_0;
(* dont_touch="true" *) wire                             l1_prio_match_0;
(* dont_touch="true" *) wire                             l1_prio_match_en_0;
assign l1_prio_match_en_0 = match_0  | match_1 ;

(* keep_hierarchy="yes" *) prio_enc1 #(
	.DATA_WIDTH (TCAM_MATCH_ADDR_WIDTH+ID_BITS)
) u_prio_enc_l1_0 (
	.clk        (clk),
	.rst_n      (rst_vct[2]),
	.en         (l1_prio_match_en_0),

	.en_0       (match_0),
	.din_0      ({match_addr_0, 1'b0}),
	.en_1       (match_1),
	.din_1      ({match_addr_1, 1'b1}),

	.dout_en    (l1_prio_match_0),
	.dout       (l1_prio_match_addr_0)
);

assign match = l1_prio_match_0;
assign match_addr = l1_prio_match_addr_0;

endmodule


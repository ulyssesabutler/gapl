module ones_complement_addition
#(
    parameter WIDTH = 16
)
(
    input  [WIDTH - 1:0] operand_1,
    input  [WIDTH - 1:0] operand_2,
    output [WIDTH - 1:0] sum
);

    // TODO

endmodule
module high_throughput_stateful_processor
#(
    parameter REPLICATION_FACTOR = 3
) (
    input  wire clock,
    input  wire reset,
    input  wire enable,

    input  wire [8 * REPLICATION_FACTOR - 1:0] data_in,
    output wire [7:0]                          data_out
);

    state_transition_main main
    (
        .clock(clock),
        .reset(reset),
        .enable(enable),

        .i(data_in),
        .o(data_out)
    );

endmodule
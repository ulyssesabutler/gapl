module one_hot_to_count
#(
    parameter INPUT_SIZE  = 32,
    localparam INDEX_BITS = $clog2(INPUT_SIZE + 2),

    localparam NEAREST_POW_2 = 2**$clog2(INPUT_SIZE)
)
(
    input      [INPUT_SIZE - 1:0] one_hot,
    output reg [INDEX_BITS - 1:0] count // Basically, one indexing
);
/*
    wire [INDEX_BITS - 1:0] bit_index;

    wire [NEAREST_POW_2 - 1:0] bit_table [INDEX_BITS - 1:0];

    genvar i;
    generate
        for (i = 0; i < INDEX_BITS; i = i + 1) begin
            assign bit_table[i] = {(NEAREST_POW_2 >> (i + 1)){{(1 << i){1'b0}}, {(1 << i){1'b1}}}};
            assign bit_index[i] = (one_hot & bit_table[i]) ? 1 : 0;
        end
    endgenerate

    assign count = one_hot ? (INPUT_SIZE - bit_index) : 0;
*/

    always @(*) begin
        case (one_hot)
            32'b00000000000000000000000000000001: count = 1;
            32'b00000000000000000000000000000010: count = 2;
            32'b00000000000000000000000000000100: count = 3;
            32'b00000000000000000000000000001000: count = 4;
            32'b00000000000000000000000000010000: count = 5;
            32'b00000000000000000000000000100000: count = 6;
            32'b00000000000000000000000001000000: count = 7;
            32'b00000000000000000000000010000000: count = 8;
            32'b00000000000000000000000100000000: count = 9;
            32'b00000000000000000000001000000000: count = 10;
            32'b00000000000000000000010000000000: count = 11;
            32'b00000000000000000000100000000000: count = 12;
            32'b00000000000000000001000000000000: count = 13;
            32'b00000000000000000010000000000000: count = 14;
            32'b00000000000000000100000000000000: count = 15;
            32'b00000000000000001000000000000000: count = 16;
            32'b00000000000000010000000000000000: count = 17;
            32'b00000000000000100000000000000000: count = 18;
            32'b00000000000001000000000000000000: count = 19;
            32'b00000000000010000000000000000000: count = 20;
            32'b00000000000100000000000000000000: count = 21;
            32'b00000000001000000000000000000000: count = 22;
            32'b00000000010000000000000000000000: count = 23;
            32'b00000000100000000000000000000000: count = 24;
            32'b00000001000000000000000000000000: count = 25;
            32'b00000010000000000000000000000000: count = 26;
            32'b00000100000000000000000000000000: count = 27;
            32'b00001000000000000000000000000000: count = 28;
            32'b00010000000000000000000000000000: count = 29;
            32'b00100000000000000000000000000000: count = 30;
            32'b01000000000000000000000000000000: count = 31;
            32'b10000000000000000000000000000000: count = 32;
            default:                              count = 0;
        endcase
    end

endmodule
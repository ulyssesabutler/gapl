//
// Copyright (C) 2019 Yuta Tokusashi
// All rights reserved.
//
// This software was developed by
// Stanford University and the University of Cambridge Computer Laboratory
// under National Science Foundation under Grant No. CNS-0855268,
// the University of Cambridge Computer Laboratory under EPSRC INTERNET Project EP/H040536/1 and
// by the University of Cambridge Computer Laboratory under DARPA/AFRL contract FA8750-11-C-0249 ("MRC2"), 
// as part of the DARPA MRC research programme.
//
// @NETFPGA_LICENSE_HEADER_START@
//
// Licensed to NetFPGA C.I.C. (NetFPGA) under one or more contributor
// license agreements.  See the NOTICE file distributed with this work for
// additional information regarding copyright ownership.  NetFPGA licenses this
// file to you under the NetFPGA Hardware-Software License, Version 1.0 (the
// "License"); you may not use this file except in compliance with the
// License.  You may obtain a copy of the License at:
//
//   http://www.netfpga-cic.org
//
// Unless required by applicable law or agreed to in writing, Work distributed
// under the License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied.  See the License for the
// specific language governing permissions and limitations under the License.
//
// @NETFPGA_LICENSE_HEADER_END@
//
 
 // This file is generated by ./gen.sh
module prio_enc1 #(
	parameter DATA_WIDTH = 32
)(
	input wire clk,
	input wire rst_n,
	input wire en,

	input wire en_0,
	input wire [DATA_WIDTH-1:0] din_0,

	input wire en_1,
	input wire [DATA_WIDTH-1:0] din_1,


	output wire                  dout_en,
	output wire [DATA_WIDTH-1:0] dout
);

 assign dout = 	(!en ) ? 0  : (
				(en_0) ? din_0 :
				(en_1) ? din_1 :
 				0);

assign dout_en = en;


endmodule

 // This file is generated by ./gen.sh
module prio_enc2 #(
	parameter DATA_WIDTH = 32
)(
	input wire clk,
	input wire rst_n,
	input wire en,

	input wire en_0,
	input wire [DATA_WIDTH-1:0] din_0,


	output wire                  dout_en,
	output wire [DATA_WIDTH-1:0] dout
);

 assign dout = 	(!en ) ? 0  : (
				(en_0) ? din_0 :
 				0);

assign dout_en = en;


endmodule

